library ieee;
use ieee.std_logic_1164.all;
use work.all;

entity uart_lcd_tester is
	port(
		
	);
end LCD_Driver;

architecture logic of LCD_Driver is